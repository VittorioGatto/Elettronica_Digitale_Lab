package State_types is
	type State_type is (A, B, C, D, E, F, G, H, I);
end State_types;