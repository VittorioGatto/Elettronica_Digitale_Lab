package State_types is
	type State_type is (A, B, C, D, E, F, G, H, I);
	type HELLO_type is (idle, start, shift1, shift2, shift3, shift4, shift5, shift6, shift7, shift8);
end State_types;