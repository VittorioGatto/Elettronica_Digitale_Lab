library ieee;
use ieee.std_logic_1164.all;
use work.serial_state_types.all;

--Behavioral implementation of look up table
entity StateLookUp is
	port(
			current_state: in State_type;
			result: out std_logic_vector(8 downto 0)
		 );
end StateLookUp;

architecture Behavior of StateLookUp is

begin
process(current_state)
begin
	case current_state is
		when A => result <= "000000001";
		when B => result <= "000000010";
		when C => result <= "000000100";
		when D => result <= "000001000";
		when E => result <= "000010000";
		when F => result <= "000100000";
		when G => result <= "001000000";
		when H => result <= "010000000";
		when I => result <= "100000000";
		when others => result <= "000000000"; --reset
	end case;
end process;
end Behavior;